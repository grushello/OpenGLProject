LevelsPassed: 4
CurrentLevel: 3
TilesTraveled: 0